/*
File containing parameters used by the modules
*/

`ifndef global_params
    `define global_params

    parameter DATA_SIZE     = 64;
    parameter ADDR_SIZE     = 32;

`endif

